-------------------------------------------------------------------------------
-- Title      : Frame checker
-- Project    : MEEP
-------------------------------------------------------------------------------
-- File        : frame_check.vhd
-- Author      : Francelly K. Cano Ladino; francelly.canoladino@bsc.es
-- Company     : Barcelona Supercomputing Center (BSC)
-- Created     : 19/01/2021 - 19:12:35
-- Last update : Mon Feb 15 13:03:35 2021
-- Synthesizer : <Name> <version>
-- FPGA        : Alveo U280
-------------------------------------------------------------------------------
-- Description:  This module will implement a Frame checker to test a loopback using Aurora 64B/66B full-duplex connection.
-- With this module, we can check the frames generated by Frame_gen that arrive from Aurora Channel (RX).
-- We used the mas pseudo data algorithm to generate the same random data as Fram_Gen, using a comparator to check both values.
-- If an error is found, there is a counter that will increment each time.
-- Signals:
--   USER_CLK: The user_clk INPUT signal is a BUFG output deriving its input from tx_out_clk (Transceivers).   
--   RESET: This INPUT  signal reset the frame checker module.
--/User Interface: RX interface
--   AXIS_UI_RX_TDATA:This input signal is the random data that come from the AXI4-stream interface
--   (Aurora Channel)
--   AXIS_UI_RX_TVALID:This input signal indicates that this modules is driving a valid transfer.
--   DATA_ERROR_COUNT:This counter indicates if the comparison was unsuccessful incrementing each time occur an unmatch.
-- Comments : <Extra comments if they were needed>
-------------------------------------------------------------------------------
-- Copyright (c) 2019 DDR/TICH
-------------------------------------------------------------------------------
-- Revisions  : 1.0
-- Date/Time                Version               Engineer
-- dd/mm/yyyy - hh:mm        1.0             francelly.canoladino@bsc.es
-- Comments   : <Highlight the modifications>
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.STD_LOGIC_1164.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;


entity frame_check is
  generic (
    DATA_WIDTH : integer := 256;
    STRB_WIDTH : integer := 32 -- STROBE bus width
    );
  port (
    -------------------------------------------------------------------------------
    -- System Interface
    -------------------------------------------------------------------------------     
    USER_CLK : in std_logic;            -- Aurora User Clk 
    RESET    : in std_logic;
    -------------------------------------------------------------------------------
    -- USER INTERFACE : RX INTERFACE
    -------------------------------------------------------------------------------
    AXIS_UI_RX_TDATA  : in  std_logic_vector(DATA_WIDTH-1 downto 0);
    AXIS_UI_RX_TVALID : in  std_logic;  --Handshake signal  
    DATA_ERR_COUNT    : out std_logic_vector(7 downto 0)
    );
end entity frame_check;

architecture rtl of frame_check is
-----------------------------------------------------------------------------
  -- CONSTANTS
-----------------------------------------------------------------------------
  constant AURORA_LANES     : integer                                      := 4;
  constant LANE_DATA_WIDTH  : integer                                      := (AURORA_LANES*64);
-----------------------------------------------------------------------------
-- SIGNALS
-----------------------------------------------------------------------------
  signal AXIS_UI_RX_TDATA_i : std_logic_vector(0 to (DATA_WIDTH-1))        := (others=>'0');
  signal r_rx_data          : std_logic_vector(0 to LANE_DATA_WIDTH-1)     := (others=>'0');
  signal r_rx_src_ready     : std_logic                                    := '0';
  signal data_err_count_r   : std_logic_vector (0 to 8-1);
  signal pdu_lfsr_r         : std_logic_vector(0 to 15)                    := (others=>'0');
  signal pdu_cmp_data_w     : std_logic_vector(LANE_DATA_WIDTH-1 downto 0) := (others=>'0');
  signal pdu_cmp_data_w_r   : std_logic_vector(0 to LANE_DATA_WIDTH-1)     := (others=>'0');
  signal data_error_c       : std_logic_vector(0 to AURORA_LANES-1)        := (others=>'0');
  signal data_error_c_r     : std_logic_vector(0 to AURORA_LANES-1)        := (others=>'0');
  signal data_error_found   : std_logic                                    := '0';
  signal data_error_not_found: std_logic                                    := '0'; 

begin

  gen_tdata : for a in 0 to STRB_WIDTH-1 generate
    AXIS_UI_RX_TDATA_i(((STRB_WIDTH-1-a)*8) to ((STRB_WIDTH-1-a)*8)+7) <= AXIS_UI_RX_TDATA(((STRB_WIDTH-1-a)*8)+7 downto ((STRB_WIDTH-1-a)*8));
  end generate gen_tdata;

  process(USER_CLK)
   begin
    if rising_edge(USER_CLK) then
      r_rx_data      <= AXIS_UI_RX_TDATA_i;
      r_rx_src_ready <= not AXIS_UI_RX_TVALID;
    end if;
  end process;
  -----------------------------------------------------------------------------
  --Pseudo data algorithm to generate the same random data as Fram_G
  ----------------------------------------------------------------------------                                      
  process(USER_CLK)
  begin
    if rising_edge(USER_CLK) then
     if RESET = '1' then
      pdu_lfsr_r <= X"ABCD";            --initial seed to start
      elsif (r_rx_src_ready = '0') then
        pdu_lfsr_r <= (not((pdu_lfsr_r(3))xor(pdu_lfsr_r(12))xor(pdu_lfsr_r(14))xor(pdu_lfsr_r(15)))&(pdu_lfsr_r(0 to 14)));
      end if;
    end if;
  end process;

  pdu_cmp_data_w <= pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&
                    pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&
                    pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&
                    pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15);
-------------------------------------------------------------------------------
-- Final data to compare
-------------------------------------------------------------------------------
  pdu_cmp_data_w_r <= pdu_cmp_data_w(255)&pdu_cmp_data_w(254)&pdu_cmp_data_w(253)&pdu_cmp_data_w(252)&
                      pdu_cmp_data_w(251)&pdu_cmp_data_w(250)&pdu_cmp_data_w(249)&pdu_cmp_data_w(248)&
                      pdu_cmp_data_w(247)&pdu_cmp_data_w(246)&pdu_cmp_data_w(245)&pdu_cmp_data_w(244)&
                      pdu_cmp_data_w(243)&pdu_cmp_data_w(242)&pdu_cmp_data_w(241)&pdu_cmp_data_w(240)&
                      pdu_cmp_data_w(239)&pdu_cmp_data_w(238)&pdu_cmp_data_w(237)&pdu_cmp_data_w(236)&
                      pdu_cmp_data_w(235)&pdu_cmp_data_w(234)&pdu_cmp_data_w(233)&pdu_cmp_data_w(232)&
                      pdu_cmp_data_w(231)&pdu_cmp_data_w(230)&pdu_cmp_data_w(229)&pdu_cmp_data_w(228)&
                      pdu_cmp_data_w(227)&pdu_cmp_data_w(226)&pdu_cmp_data_w(225)&pdu_cmp_data_w(224)&
                      pdu_cmp_data_w(223)&pdu_cmp_data_w(222)&pdu_cmp_data_w(221)&pdu_cmp_data_w(220)&
                      pdu_cmp_data_w(219)&pdu_cmp_data_w(218)&pdu_cmp_data_w(217)&pdu_cmp_data_w(216)&
                      pdu_cmp_data_w(215)&pdu_cmp_data_w(214)&pdu_cmp_data_w(213)&pdu_cmp_data_w(212)&
                      pdu_cmp_data_w(211)&pdu_cmp_data_w(210)&pdu_cmp_data_w(209)&pdu_cmp_data_w(208)&
                      pdu_cmp_data_w(207)&pdu_cmp_data_w(206)&pdu_cmp_data_w(205)&pdu_cmp_data_w(204)&
                      pdu_cmp_data_w(203)&pdu_cmp_data_w(202)&pdu_cmp_data_w(201)&pdu_cmp_data_w(200)&
                      pdu_cmp_data_w(199)&pdu_cmp_data_w(198)&pdu_cmp_data_w(197)&pdu_cmp_data_w(196)&
                      pdu_cmp_data_w(195)&pdu_cmp_data_w(194)&pdu_cmp_data_w(193)&pdu_cmp_data_w(192)&
                      pdu_cmp_data_w(191)&pdu_cmp_data_w(190)&pdu_cmp_data_w(189)&pdu_cmp_data_w(188)&--
                      pdu_cmp_data_w(187)&pdu_cmp_data_w(186)&pdu_cmp_data_w(185)&pdu_cmp_data_w(184)&
                      pdu_cmp_data_w(183)&pdu_cmp_data_w(182)&pdu_cmp_data_w(181)&pdu_cmp_data_w(180)&
                      pdu_cmp_data_w(179)&pdu_cmp_data_w(178)&pdu_cmp_data_w(177)&pdu_cmp_data_w(176)&
                      pdu_cmp_data_w(175)&pdu_cmp_data_w(174)&pdu_cmp_data_w(173)&pdu_cmp_data_w(172)&
                      pdu_cmp_data_w(171)&pdu_cmp_data_w(170)&pdu_cmp_data_w(169)&pdu_cmp_data_w(168)&
                      pdu_cmp_data_w(167)&pdu_cmp_data_w(166)&pdu_cmp_data_w(165)&pdu_cmp_data_w(164)&
                      pdu_cmp_data_w(163)&pdu_cmp_data_w(162)&pdu_cmp_data_w(161)&pdu_cmp_data_w(160)&
                      pdu_cmp_data_w(159)&pdu_cmp_data_w(158)&pdu_cmp_data_w(157)&pdu_cmp_data_w(156)&
                      pdu_cmp_data_w(155)&pdu_cmp_data_w(154)&pdu_cmp_data_w(153)&pdu_cmp_data_w(152)&
                      pdu_cmp_data_w(151)&pdu_cmp_data_w(150)&pdu_cmp_data_w(149)&pdu_cmp_data_w(148)&
                      pdu_cmp_data_w(147)&pdu_cmp_data_w(146)&pdu_cmp_data_w(145)&pdu_cmp_data_w(144)&
                      pdu_cmp_data_w(143)&pdu_cmp_data_w(142)&pdu_cmp_data_w(141)&pdu_cmp_data_w(140)&
                      pdu_cmp_data_w(139)&pdu_cmp_data_w(138)&pdu_cmp_data_w(137)&pdu_cmp_data_w(136)&
                      pdu_cmp_data_w(135)&pdu_cmp_data_w(134)&pdu_cmp_data_w(133)&pdu_cmp_data_w(132)&
                      pdu_cmp_data_w(131)&pdu_cmp_data_w(130)&pdu_cmp_data_w(129)&pdu_cmp_data_w(128)&
                      pdu_cmp_data_w(127)&pdu_cmp_data_w(126)&pdu_cmp_data_w(125)&pdu_cmp_data_w(124)&--
                      pdu_cmp_data_w(123)&pdu_cmp_data_w(122)&pdu_cmp_data_w(121)&pdu_cmp_data_w(120)&
                      pdu_cmp_data_w(119)&pdu_cmp_data_w(118)&pdu_cmp_data_w(117)&pdu_cmp_data_w(116)&
                      pdu_cmp_data_w(115)&pdu_cmp_data_w(114)&pdu_cmp_data_w(113)&pdu_cmp_data_w(112)&
                      pdu_cmp_data_w(111)&pdu_cmp_data_w(110)&pdu_cmp_data_w(109)&pdu_cmp_data_w(108)&
                      pdu_cmp_data_w(107)&pdu_cmp_data_w(106)&pdu_cmp_data_w(105)&pdu_cmp_data_w(104)&
                      pdu_cmp_data_w(103)&pdu_cmp_data_w(102)&pdu_cmp_data_w(101)&pdu_cmp_data_w(100)&
                      pdu_cmp_data_w(99)&pdu_cmp_data_w(98)&pdu_cmp_data_w(97)&pdu_cmp_data_w(96)&
                      pdu_cmp_data_w(95)&pdu_cmp_data_w(94)&pdu_cmp_data_w(93)&pdu_cmp_data_w(92)&
                      pdu_cmp_data_w(91)&pdu_cmp_data_w(90)&pdu_cmp_data_w(89)&pdu_cmp_data_w(88)&
                      pdu_cmp_data_w(87)&pdu_cmp_data_w(86)&pdu_cmp_data_w(85)&pdu_cmp_data_w(84)&
                      pdu_cmp_data_w(83)&pdu_cmp_data_w(82)&pdu_cmp_data_w(81)&pdu_cmp_data_w(80)&
                      pdu_cmp_data_w(79)&pdu_cmp_data_w(78)&pdu_cmp_data_w(77)&pdu_cmp_data_w(76)&
                      pdu_cmp_data_w(75)&pdu_cmp_data_w(74)&pdu_cmp_data_w(73)&pdu_cmp_data_w(72)&
                      pdu_cmp_data_w(71)&pdu_cmp_data_w(70)&pdu_cmp_data_w(69)&pdu_cmp_data_w(68)&
                      pdu_cmp_data_w(67)&pdu_cmp_data_w(66)&pdu_cmp_data_w(65)&pdu_cmp_data_w(64)&
                      pdu_cmp_data_w(63)&pdu_cmp_data_w(62)&pdu_cmp_data_w(61)&pdu_cmp_data_w(60)&--
                      pdu_cmp_data_w(59)&pdu_cmp_data_w(58)&pdu_cmp_data_w(57)&pdu_cmp_data_w(56)&
                      pdu_cmp_data_w(55)&pdu_cmp_data_w(54)&pdu_cmp_data_w(53)&pdu_cmp_data_w(52)&
                      pdu_cmp_data_w(51)&pdu_cmp_data_w(50)&pdu_cmp_data_w(49)&pdu_cmp_data_w(48)&
                      pdu_cmp_data_w(47)&pdu_cmp_data_w(46)&pdu_cmp_data_w(45)&pdu_cmp_data_w(44)&
                      pdu_cmp_data_w(43)&pdu_cmp_data_w(42)&pdu_cmp_data_w(41)&pdu_cmp_data_w(40)&
                      pdu_cmp_data_w(39)&pdu_cmp_data_w(38)&pdu_cmp_data_w(37)&pdu_cmp_data_w(36)&
                      pdu_cmp_data_w(35)&pdu_cmp_data_w(34)&pdu_cmp_data_w(33)&pdu_cmp_data_w(32)&
                      pdu_cmp_data_w(31)&pdu_cmp_data_w(30)&pdu_cmp_data_w(29)&pdu_cmp_data_w(28)&
                      pdu_cmp_data_w(27)&pdu_cmp_data_w(26)&pdu_cmp_data_w(25)&pdu_cmp_data_w(24)&
                      pdu_cmp_data_w(23)&pdu_cmp_data_w(22)&pdu_cmp_data_w(21)&pdu_cmp_data_w(20)&
                      pdu_cmp_data_w(19)&pdu_cmp_data_w(18)&pdu_cmp_data_w(17)&pdu_cmp_data_w(16)&
                      pdu_cmp_data_w(15)&pdu_cmp_data_w(14)&pdu_cmp_data_w(13)&pdu_cmp_data_w(12)&
                      pdu_cmp_data_w(11)&pdu_cmp_data_w(10)&pdu_cmp_data_w(9)&pdu_cmp_data_w(8)&
                      pdu_cmp_data_w(7)&pdu_cmp_data_w(6)&pdu_cmp_data_w(5)&pdu_cmp_data_w(4)&
                      pdu_cmp_data_w(3)&pdu_cmp_data_w(2)&pdu_cmp_data_w(1)&pdu_cmp_data_w(0);
-- Data error counter

data_error_c(0)<='1' when ( (r_rx_src_ready='0') and (r_rx_data(0 to 63)/=pdu_cmp_data_w_r(0 to 63))) else
                 '0';
             
process(USER_CLK)
 begin
   if rising_edge(USER_CLK) then  
     data_error_c_r<=  data_error_c;    
end if;
end process;

data_error_not_found<=data_err_count_r(0) and data_err_count_r(1) and data_err_count_r(2) and data_err_count_r(3) and data_err_count_r(4) and data_err_count_r(5) and data_err_count_r(6) and data_err_count_r(7);
--data_error_found<=data_error_c_r(3) or data_error_c_r(2) or data_error_c_r(1) or data_error_c_r(0);-- or data_err_c_r(4) or data_err_c_r(5) or data_err_c_r(6) or data_err_c_r(7);
data_error_found<=data_error_c(0);-- or data_error_c_r(2) or data_error_c_r(1) or data_error_c_r(0);

process(USER_CLK)
 begin
   if rising_edge(USER_CLK) then
	 if RESET ='1' then
		data_err_count_r <=(others=> '0'); 
	   elsif data_err_count_r= 255  then
	      --data_err_count_r<=data_err_count_r;	
	      data_err_count_r <=(others=> '0');     
		elsif data_error_found ='1' then
			data_err_count_r <= data_err_count_r + 1;
		end if;
   end if;
end process;

--process(USER_CLK)
--begin
--	if rising_edge(USER_CLK) then
--	 if RESET ='1' then
--		data_err_count_r <=(others=> '0'); 
--	   elsif r_rx_src_ready='0' then
--	    if  data_err_count_r= 255 then
--	       data_err_count_r <=(others=> '0'); 
--		elsif (pdu_cmp_data_w_r/=r_rx_data ) then
--			data_err_count_r <= data_err_count_r + 1;
--		end if;
--	end if; 
--end if;
--end process;

DATA_ERR_COUNT<=data_err_count_r;

end architecture rtl;
